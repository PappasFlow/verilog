`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:33:00 08/23/2022 
// Design Name: 
// Module Name:    Act4_VM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Act4_VM(
    input A,
    input B,
    input C,
    output F1,
    output F2,
    output F3,
    output F4
    );


and (F1,~A,B);


endmodule
